module Contador (
    input  wire clk,
    input  wire rst_n,

    input  wire acrescer,
    input  wire decrecer,

    output wire [7:0] saida
);

// Insira seu código aqui

endmodule
